module adder(input []data1, data2  ,output bpc);
	assign bpc = data1+data2;
endmodule
