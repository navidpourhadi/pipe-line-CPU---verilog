module adder(input [63:0]data1 , data2  ,output[63:0] result);
	assign result = data1+data2;
endmodule
