module adder(input apc  ,output bpc);
	assign bpc = apc+4;
endmodule
